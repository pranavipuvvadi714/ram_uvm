`include "interface.sv"
`include "ram_defines.svh"
package ram_pkg;
`include "ram_trans.sv"
`include "ram_wr_seq.sv"
`include "ram_rd_seq.sv"
`include "ram_wr_sequencer.sv"
`include "ram_rd_sequencer.sv"
`include "ram_wr_driver.sv"
`include "ram_rd_driver.sv"
`include "ram_wr_monitor.sv"
`include "ram_rd_monitor.sv"
`include "ram_wr_agent.sv"
`include "ram_rd_agent.sv"
`include "ram_env.sv"
`include "ram_scoreboard.sv"
`include "ram_base_test.sv"
endpackage
