`define ADDR_WIDTH 4
`define DATA_WIDTH 8
`define DEPTH 16
`define no_of_itr 20
